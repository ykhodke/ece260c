package utopia_pkg;
  `import uvm_pkg::*;
  `include "uvm_macros.svh"

  `define TxPorts 4 //set number of transmit ports
  `define RxPorts 4 //set number of receive ports

  parameter NumTx = `TxPorts;
  parameter NumRx = `RxPorts;


/* ## Cell definition formats go here ## */
  
  /* UNI cell format */
  typedef struct packed {
    bit        [3:0]  GFC;
    bit        [7:0]  VPI;
    bit        [15:0] VCI;
    bit               CLP;
    bit        [2:0]  PT;
    bit        [7:0]  HEC;
    bit [0:47] [7:0]  Payload;
  } uniType;

  /* NNI Cell Format */
  typedef struct packed {
    bit        [11:0] VPI;
    bit        [15:0] VCI;
    bit               CLP;
    bit        [2:0]  PT;
    bit        [7:0]  HEC;
    bit [0:47] [7:0]  Payload;
  } nniType;

  /* Test View Cell Format (Payload Section) */
  typedef struct packed {
    bit [0:4]  [7:0] Header;
    bit [0:3]  [7:0] PortID;
    bit [0:3]  [7:0] CellID;
    bit [0:39] [7:0] Padding;
  } tstType;

  /* Union of UNI / NNI / Test View / ByteStream */
  typedef union packed {
    uniType uni;
    nniType nni;
    tstType tst;
    bit [0:52] [7:0] Mem;
  } ATMCellType;

  /* Cell Rewriting and Forwarding Configuration */
  typedef struct packed {
    bit [`TxPorts-1:0] FWD;
    bit [11:0] VPI;
  } CellCfgType;



/* ## included header files go here ## */

  `include "coverage.svh"
  `include "scoreboard.svh"

  // TODO :: include the rest of the moduel definitions here 


endpackage : utopia_pkg